module vxlsx_io

#flag -lxlsxio_read
#include <xlsxio_read.h>

#flag -lxlsxio_write
#include <xlsxio_write.h>

pub const vxlsx_io_null = unsafe { nil }
