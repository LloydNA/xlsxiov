module vxlsxio

#flag -lxlsxio_read
#include <xlsxio_read.h>

#flag -lxlsxio_write
#include <xlsxio_write.h>

pub const vxlsxio_null = unsafe { nil }
